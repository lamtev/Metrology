** Profile: "SCHEMATIC1-watts"  [ D:\metrology\power_regulator\orcad\modeling_schema\schema-schematic1-watts.sim ] 

** Creating circuit file "schema-schematic1-watts.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.STMLIB ".\SCHEMA.stl" 
* From [PSPICE NETLIST] section of C:\Programs\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 20ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\schema-SCHEMATIC1.net" 


.END
