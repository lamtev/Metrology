** Profile: "SCHEMATIC1-220sin50"  [ D:\METROLOGY\POWER_REGULATOR\ORCAD\pow_reg-SCHEMATIC1-220sin50.sim ] 

** Creating circuit file "pow_reg-SCHEMATIC1-220sin50.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.STMLIB ".\POW_REG.stl" 
* From [PSPICE NETLIST] section of C:\Programs\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 60ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\pow_reg-SCHEMATIC1.net" 


.END
