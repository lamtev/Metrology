** Profile: "SCHEMATIC1-rect_imp"  [ D:\metrology\rc_int_circuit\rc_int_circuit-schematic1-rect_imp.sim ] 

** Creating circuit file "rc_int_circuit-schematic1-rect_imp.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
.STMLIB ".\RC_INT_CIRCUIT.stl" 
* From [PSPICE NETLIST] section of C:\Programs\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 3u 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\rc_int_circuit-SCHEMATIC1.net" 


.END
